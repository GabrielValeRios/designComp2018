-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 17.1.0 Build 590 10/25/2017 SJ Lite Edition
-- Created on Thu Oct 04 21:52:59 2018

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SMUC IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        Z : IN STD_LOGIC := '0';
        ft : IN STD_LOGIC := '0';
        iniciaMaquina : IN STD_LOGIC := '0';
        resets : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
        enables : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
        SelULA : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        SelMUX : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        number : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END SMUC;

ARCHITECTURE BEHAVIOR OF SMUC IS
    TYPE type_fstate IS (us,ds,um,dm,uh,dh,UsDs10,DsUm6,UmDm10,DmUh6,UhDh10,waitState);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_resets : STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
    SIGNAL reg_enables : STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
    SIGNAL reg_SelULA : STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
    SIGNAL reg_SelMUX : STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
    SIGNAL reg_number : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Z,ft,iniciaMaquina,reg_resets,reg_enables,reg_SelULA,reg_SelMUX,reg_number)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= waitState;
            reg_resets <= "000000";
            reg_enables <= "000000";
            reg_SelULA <= "000";
            reg_SelMUX <= "000";
            reg_number <= "0000";
            resets <= "000000";
            enables <= "000000";
            SelULA <= "000";
            SelMUX <= "000";
            number <= "0000";
        ELSE
            reg_resets <= "000000";
            reg_enables <= "000000";
            reg_SelULA <= "000";
            reg_SelMUX <= "000";
            reg_number <= "0000";
            resets <= "000000";
            enables <= "000000";
            SelULA <= "000";
            SelMUX <= "000";
            number <= "0000";
            CASE fstate IS
                WHEN us =>
                    IF ((ft = '1')) THEN
                        reg_fstate <= UsDs10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= us;
                    END IF;

                    reg_SelULA <= "001";

                    reg_SelMUX <= "000";

                    reg_enables <= "000001";

                    reg_resets <= "000000";

                    reg_number <= "0001";
                WHEN ds =>
                    IF ((ft = '1')) THEN
                        reg_fstate <= DsUm6;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ds;
                    END IF;

                    reg_SelULA <= "001";

                    reg_SelMUX <= "001";

                    reg_enables <= "000010";

                    reg_resets <= "000001";

                    reg_number <= "0001";
                WHEN um =>
                    IF ((ft = '1')) THEN
                        reg_fstate <= UmDm10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= um;
                    END IF;

                    reg_SelULA <= "001";

                    reg_SelMUX <= "010";

                    reg_enables <= "000100";

                    reg_resets <= "000011";

                    reg_number <= "0001";
                WHEN dm =>
                    IF ((ft = '1')) THEN
                        reg_fstate <= DmUh6;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= dm;
                    END IF;

                    reg_SelULA <= "001";

                    reg_SelMUX <= "011";

                    reg_enables <= "001000";

                    reg_resets <= "000111";

                    reg_number <= "0001";
                WHEN uh =>
                    IF ((ft = '1')) THEN
                        reg_fstate <= UhDh10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= uh;
                    END IF;

                    reg_SelULA <= "001";

                    reg_SelMUX <= "100";

                    reg_enables <= "010000";

                    reg_resets <= "001111";

                    reg_number <= "0001";
                WHEN dh =>
                    IF ((ft = '1')) THEN
                        reg_fstate <= waitState;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= dh;
                    END IF;

                    reg_SelULA <= "001";

                    reg_SelMUX <= "101";

                    reg_enables <= "100000";

                    reg_resets <= "011111";

                    reg_number <= "0001";
                WHEN UsDs10 =>
                    IF (NOT((Z = '1'))) THEN
                        reg_fstate <= waitState;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= ds;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= UsDs10;
                    END IF;

                    reg_SelULA <= "010";

                    reg_SelMUX <= "000";

                    reg_number <= "1010";
                WHEN DsUm6 =>
                    IF (NOT((Z = '1'))) THEN
                        reg_fstate <= waitState;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= um;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= DsUm6;
                    END IF;

                    reg_SelULA <= "010";

                    reg_SelMUX <= "001";

                    reg_number <= "0110";
                WHEN UmDm10 =>
                    IF (NOT((Z = '1'))) THEN
                        reg_fstate <= waitState;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= dm;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= UmDm10;
                    END IF;

                    reg_SelULA <= "010";

                    reg_SelMUX <= "010";

                    reg_number <= "1010";
                WHEN DmUh6 =>
                    IF (NOT((Z = '1'))) THEN
                        reg_fstate <= waitState;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= uh;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= DmUh6;
                    END IF;

                    reg_SelULA <= "010";

                    reg_SelMUX <= "011";

                    reg_number <= "0110";
                WHEN UhDh10 =>
                    IF (NOT((Z = '1'))) THEN
                        reg_fstate <= waitState;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= dh;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= UhDh10;
                    END IF;

                    reg_SelULA <= "010";

                    reg_SelMUX <= "100";

                    reg_number <= "1010";
                WHEN waitState =>
                    IF (NOT((iniciaMaquina = '1'))) THEN
                        reg_fstate <= waitState;
                    ELSIF ((iniciaMaquina = '1')) THEN
                        reg_fstate <= us;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= waitState;
                    END IF;

                    reg_number <= "0000";
                WHEN OTHERS => 
                    reg_resets <= "XXXXXX";
                    reg_enables <= "XXXXXX";
                    reg_SelULA <= "XXX";
                    reg_SelMUX <= "XXX";
                    reg_number <= "XXXX";
                    report "Reach undefined state";
            END CASE;
            resets <= reg_resets;
            enables <= reg_enables;
            SelULA <= reg_SelULA;
            SelMUX <= reg_SelMUX;
            number <= reg_number;
        END IF;
    END PROCESS;
END BEHAVIOR;
