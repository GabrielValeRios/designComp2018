-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Intel and sold by Intel or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 17.0.0 Build 595 04/25/2017 SJ Lite Edition
-- Created on Tue Oct 10 21:25:10 2017

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SM IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        bt1 : IN STD_LOGIC := '0';
        bt2 : IN STD_LOGIC := '0';
        bt3 : IN STD_LOGIC := '0';
        saida : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
END SM;

ARCHITECTURE BEHAVIOR OF SM IS
    TYPE type_fstate IS (state0,state1,state2);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_saida : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,bt1,bt2,bt3,reg_saida)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state0;
            reg_saida <= "0000";
            saida <= "0000";
        ELSE
            reg_saida <= "0000";
            saida <= "0000";
            CASE fstate IS
                WHEN state0 =>
                    IF (((NOT((bt1 = '1')) AND (bt2 = '1')) AND NOT((bt3 = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF (((NOT((bt1 = '1')) AND NOT((bt2 = '1'))) AND (bt3 = '1'))) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state0;
                    END IF;

                    reg_saida <= "0000";
                WHEN state1 =>
                    IF (((NOT((bt1 = '1')) AND NOT((bt2 = '1'))) AND (bt3 = '1'))) THEN
                        reg_fstate <= state2;
                    ELSIF ((((bt1 = '1') AND NOT((bt2 = '1'))) AND NOT((bt3 = '1')))) THEN
                        reg_fstate <= state0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    reg_saida <= "0001";
                WHEN state2 =>
                    IF (((NOT((bt1 = '1')) AND (bt2 = '1')) AND NOT((bt3 = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF ((((bt1 = '1') AND NOT((bt2 = '1'))) AND NOT((bt3 = '1')))) THEN
                        reg_fstate <= state0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    reg_saida <= "0010";
                WHEN OTHERS => 
                    reg_saida <= "XXXX";
                    report "Reach undefined state";
            END CASE;
            saida <= reg_saida;
        END IF;
    END PROCESS;
END BEHAVIOR;
